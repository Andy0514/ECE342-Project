
module PROBE_1 (
	source,
	probe,
	source_clk);	

	output	[0:0]	source;
	input	[0:0]	probe;
	input		source_clk;
endmodule
