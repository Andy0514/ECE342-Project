
module PROBE_32 (
	probe);	

	input	[31:0]	probe;
endmodule
