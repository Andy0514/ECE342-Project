
module PROBE_256 (
	source,
	source_clk);	

	output	[255:0]	source;
	input		source_clk;
endmodule
