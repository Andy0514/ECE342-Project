
module PROBE_96 (
	source,
	source_clk);	

	output	[95:0]	source;
	input		source_clk;
endmodule
